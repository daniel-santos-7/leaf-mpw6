magic
tech sky130A
magscale 1 2
timestamp 1652032400
<< nwell >>
rect 1066 276613 278890 277179
rect 1066 275525 278890 276091
rect 1066 274437 278890 275003
rect 1066 273349 278890 273915
rect 1066 272261 278890 272827
rect 1066 271173 278890 271739
rect 1066 270085 278890 270651
rect 1066 268997 278890 269563
rect 1066 267909 278890 268475
rect 1066 266821 278890 267387
rect 1066 265733 278890 266299
rect 1066 264645 278890 265211
rect 1066 263557 278890 264123
rect 1066 262469 278890 263035
rect 1066 261381 278890 261947
rect 1066 260293 278890 260859
rect 1066 259205 278890 259771
rect 1066 258117 278890 258683
rect 1066 257029 278890 257595
rect 1066 255941 278890 256507
rect 1066 254853 278890 255419
rect 1066 253765 278890 254331
rect 1066 252677 278890 253243
rect 1066 251589 278890 252155
rect 1066 250501 278890 251067
rect 1066 249413 278890 249979
rect 1066 248325 278890 248891
rect 1066 247237 278890 247803
rect 1066 246149 278890 246715
rect 1066 245061 278890 245627
rect 1066 243973 278890 244539
rect 1066 242885 278890 243451
rect 1066 241797 278890 242363
rect 1066 240709 278890 241275
rect 1066 239621 278890 240187
rect 1066 238533 278890 239099
rect 1066 237445 278890 238011
rect 1066 236357 278890 236923
rect 1066 235269 278890 235835
rect 1066 234181 278890 234747
rect 1066 233093 278890 233659
rect 1066 232005 278890 232571
rect 1066 230917 278890 231483
rect 1066 229829 278890 230395
rect 1066 228741 278890 229307
rect 1066 227653 278890 228219
rect 1066 226565 278890 227131
rect 1066 225477 278890 226043
rect 1066 224389 278890 224955
rect 1066 223301 278890 223867
rect 1066 222213 278890 222779
rect 1066 221125 278890 221691
rect 1066 220037 278890 220603
rect 1066 218949 278890 219515
rect 1066 217861 278890 218427
rect 1066 216773 278890 217339
rect 1066 215685 278890 216251
rect 1066 214597 278890 215163
rect 1066 213509 278890 214075
rect 1066 212421 278890 212987
rect 1066 211333 278890 211899
rect 1066 210245 278890 210811
rect 1066 209157 278890 209723
rect 1066 208069 278890 208635
rect 1066 206981 278890 207547
rect 1066 205893 278890 206459
rect 1066 204805 278890 205371
rect 1066 203717 278890 204283
rect 1066 202629 278890 203195
rect 1066 201541 278890 202107
rect 1066 200453 278890 201019
rect 1066 199365 278890 199931
rect 1066 198277 278890 198843
rect 1066 197189 278890 197755
rect 1066 196101 278890 196667
rect 1066 195013 278890 195579
rect 1066 193925 278890 194491
rect 1066 192837 278890 193403
rect 1066 191749 278890 192315
rect 1066 190661 278890 191227
rect 1066 189573 278890 190139
rect 1066 188485 278890 189051
rect 1066 187397 278890 187963
rect 1066 186309 278890 186875
rect 1066 185221 278890 185787
rect 1066 184133 278890 184699
rect 1066 183045 278890 183611
rect 1066 181957 278890 182523
rect 1066 180869 278890 181435
rect 1066 179781 278890 180347
rect 1066 178693 278890 179259
rect 1066 177605 278890 178171
rect 1066 176517 278890 177083
rect 1066 175429 278890 175995
rect 1066 174341 278890 174907
rect 1066 173253 278890 173819
rect 1066 172165 278890 172731
rect 1066 171077 278890 171643
rect 1066 169989 278890 170555
rect 1066 168901 278890 169467
rect 1066 167813 278890 168379
rect 1066 166725 278890 167291
rect 1066 165637 278890 166203
rect 1066 164549 278890 165115
rect 1066 163461 278890 164027
rect 1066 162373 278890 162939
rect 1066 161285 278890 161851
rect 1066 160197 278890 160763
rect 1066 159109 278890 159675
rect 1066 158021 278890 158587
rect 1066 156933 278890 157499
rect 1066 155845 278890 156411
rect 1066 154757 278890 155323
rect 1066 153669 278890 154235
rect 1066 152581 278890 153147
rect 1066 151493 278890 152059
rect 1066 150405 278890 150971
rect 1066 149317 278890 149883
rect 1066 148229 278890 148795
rect 1066 147141 278890 147707
rect 1066 146053 278890 146619
rect 1066 144965 278890 145531
rect 1066 143877 278890 144443
rect 1066 142789 278890 143355
rect 1066 141701 278890 142267
rect 1066 140613 278890 141179
rect 1066 139525 278890 140091
rect 1066 138437 278890 139003
rect 1066 137349 278890 137915
rect 1066 136261 278890 136827
rect 1066 135173 278890 135739
rect 1066 134085 278890 134651
rect 1066 132997 278890 133563
rect 1066 131909 278890 132475
rect 1066 130821 278890 131387
rect 1066 129733 278890 130299
rect 1066 128645 278890 129211
rect 1066 127557 278890 128123
rect 1066 126469 278890 127035
rect 1066 125381 278890 125947
rect 1066 124293 278890 124859
rect 1066 123205 278890 123771
rect 1066 122117 278890 122683
rect 1066 121029 278890 121595
rect 1066 119941 278890 120507
rect 1066 118853 278890 119419
rect 1066 117765 278890 118331
rect 1066 116677 278890 117243
rect 1066 115589 278890 116155
rect 1066 114501 278890 115067
rect 1066 113413 278890 113979
rect 1066 112325 278890 112891
rect 1066 111237 278890 111803
rect 1066 110149 278890 110715
rect 1066 109061 278890 109627
rect 1066 107973 278890 108539
rect 1066 106885 278890 107451
rect 1066 105797 278890 106363
rect 1066 104709 278890 105275
rect 1066 103621 278890 104187
rect 1066 102533 278890 103099
rect 1066 101445 278890 102011
rect 1066 100357 278890 100923
rect 1066 99269 278890 99835
rect 1066 98181 278890 98747
rect 1066 97093 278890 97659
rect 1066 96005 278890 96571
rect 1066 94917 278890 95483
rect 1066 93829 278890 94395
rect 1066 92741 278890 93307
rect 1066 91653 278890 92219
rect 1066 90565 278890 91131
rect 1066 89477 278890 90043
rect 1066 88389 278890 88955
rect 1066 87301 278890 87867
rect 1066 86213 278890 86779
rect 1066 85125 278890 85691
rect 1066 84037 278890 84603
rect 1066 82949 278890 83515
rect 1066 81861 278890 82427
rect 1066 80773 278890 81339
rect 1066 79685 278890 80251
rect 1066 78597 278890 79163
rect 1066 77509 278890 78075
rect 1066 76421 278890 76987
rect 1066 75333 278890 75899
rect 1066 74245 278890 74811
rect 1066 73157 278890 73723
rect 1066 72069 278890 72635
rect 1066 70981 278890 71547
rect 1066 69893 278890 70459
rect 1066 68805 278890 69371
rect 1066 67717 278890 68283
rect 1066 66629 278890 67195
rect 1066 65541 278890 66107
rect 1066 64453 278890 65019
rect 1066 63365 278890 63931
rect 1066 62277 278890 62843
rect 1066 61189 278890 61755
rect 1066 60101 278890 60667
rect 1066 59013 278890 59579
rect 1066 57925 278890 58491
rect 1066 56837 278890 57403
rect 1066 55749 278890 56315
rect 1066 54661 278890 55227
rect 1066 53573 278890 54139
rect 1066 52485 278890 53051
rect 1066 51397 278890 51963
rect 1066 50309 278890 50875
rect 1066 49221 278890 49787
rect 1066 48133 278890 48699
rect 1066 47045 278890 47611
rect 1066 45957 278890 46523
rect 1066 44869 278890 45435
rect 1066 43781 278890 44347
rect 1066 42693 278890 43259
rect 1066 41605 278890 42171
rect 1066 40517 278890 41083
rect 1066 39429 278890 39995
rect 1066 38341 278890 38907
rect 1066 37253 278890 37819
rect 1066 36165 278890 36731
rect 1066 35077 278890 35643
rect 1066 33989 278890 34555
rect 1066 32901 278890 33467
rect 1066 31813 278890 32379
rect 1066 30725 278890 31291
rect 1066 29637 278890 30203
rect 1066 28549 278890 29115
rect 1066 27461 278890 28027
rect 1066 26373 278890 26939
rect 1066 25285 278890 25851
rect 1066 24197 278890 24763
rect 1066 23109 278890 23675
rect 1066 22021 278890 22587
rect 1066 20933 278890 21499
rect 1066 19845 278890 20411
rect 1066 18757 278890 19323
rect 1066 17669 278890 18235
rect 1066 16581 278890 17147
rect 1066 15493 278890 16059
rect 1066 14405 278890 14971
rect 1066 13317 278890 13883
rect 1066 12229 278890 12795
rect 1066 11141 278890 11707
rect 1066 10053 278890 10619
rect 1066 8965 278890 9531
rect 1066 7877 278890 8443
rect 1066 6789 278890 7355
rect 1066 5701 278890 6267
rect 1066 4613 278890 5179
rect 1066 3525 278890 4091
rect 1066 2437 278890 3003
<< obsli1 >>
rect 1104 2159 278852 277457
<< obsm1 >>
rect 1104 2128 278852 277488
<< metal2 >>
rect 69938 279200 69994 280000
rect 209870 279200 209926 280000
rect 69938 0 69994 800
rect 209870 0 209926 800
<< obsm2 >>
rect 1860 279144 69882 279200
rect 70050 279144 209814 279200
rect 209982 279144 278004 279200
rect 1860 856 278004 279144
rect 1860 800 69882 856
rect 70050 800 209814 856
rect 209982 800 278004 856
<< obsm3 >>
rect 2957 2143 276999 277473
<< metal4 >>
rect 4208 2128 4528 277488
rect 19568 2128 19888 277488
rect 34928 2128 35248 277488
rect 50288 2128 50608 277488
rect 65648 2128 65968 277488
rect 81008 2128 81328 277488
rect 96368 2128 96688 277488
rect 111728 2128 112048 277488
rect 127088 2128 127408 277488
rect 142448 2128 142768 277488
rect 157808 2128 158128 277488
rect 173168 2128 173488 277488
rect 188528 2128 188848 277488
rect 203888 2128 204208 277488
rect 219248 2128 219568 277488
rect 234608 2128 234928 277488
rect 249968 2128 250288 277488
rect 265328 2128 265648 277488
<< obsm4 >>
rect 18827 2347 19488 265573
rect 19968 2347 34848 265573
rect 35328 2347 50208 265573
rect 50688 2347 65568 265573
rect 66048 2347 80928 265573
rect 81408 2347 96288 265573
rect 96768 2347 111648 265573
rect 112128 2347 127008 265573
rect 127488 2347 142368 265573
rect 142848 2347 157728 265573
rect 158208 2347 173088 265573
rect 173568 2347 188448 265573
rect 188928 2347 203808 265573
rect 204288 2347 219168 265573
rect 219648 2347 234528 265573
rect 235008 2347 249888 265573
rect 250368 2347 265248 265573
rect 265728 2347 275757 265573
<< labels >>
rlabel metal2 s 69938 0 69994 800 6 clk
port 1 nsew signal input
rlabel metal2 s 209870 0 209926 800 6 reset
port 2 nsew signal input
rlabel metal2 s 69938 279200 69994 280000 6 rx
port 3 nsew signal input
rlabel metal2 s 209870 279200 209926 280000 6 tx
port 4 nsew signal output
rlabel metal4 s 4208 2128 4528 277488 6 vccd1
port 5 nsew power input
rlabel metal4 s 34928 2128 35248 277488 6 vccd1
port 5 nsew power input
rlabel metal4 s 65648 2128 65968 277488 6 vccd1
port 5 nsew power input
rlabel metal4 s 96368 2128 96688 277488 6 vccd1
port 5 nsew power input
rlabel metal4 s 127088 2128 127408 277488 6 vccd1
port 5 nsew power input
rlabel metal4 s 157808 2128 158128 277488 6 vccd1
port 5 nsew power input
rlabel metal4 s 188528 2128 188848 277488 6 vccd1
port 5 nsew power input
rlabel metal4 s 219248 2128 219568 277488 6 vccd1
port 5 nsew power input
rlabel metal4 s 249968 2128 250288 277488 6 vccd1
port 5 nsew power input
rlabel metal4 s 19568 2128 19888 277488 6 vssd1
port 6 nsew ground input
rlabel metal4 s 50288 2128 50608 277488 6 vssd1
port 6 nsew ground input
rlabel metal4 s 81008 2128 81328 277488 6 vssd1
port 6 nsew ground input
rlabel metal4 s 111728 2128 112048 277488 6 vssd1
port 6 nsew ground input
rlabel metal4 s 142448 2128 142768 277488 6 vssd1
port 6 nsew ground input
rlabel metal4 s 173168 2128 173488 277488 6 vssd1
port 6 nsew ground input
rlabel metal4 s 203888 2128 204208 277488 6 vssd1
port 6 nsew ground input
rlabel metal4 s 234608 2128 234928 277488 6 vssd1
port 6 nsew ground input
rlabel metal4 s 265328 2128 265648 277488 6 vssd1
port 6 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 280000 280000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 99902758
string GDS_FILE /home/daniel-lx/caravel-mpw-6b/mpw-6b/openlane/leaf_chip/runs/leaf_chip/results/finishing/leaf_chip.magic.gds
string GDS_START 1678128
<< end >>

