VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO leaf_chip
  CLASS BLOCK ;
  FOREIGN leaf_chip ;
  ORIGIN 0.000 0.000 ;
  SIZE 1400.000 BY 1400.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 349.690 0.000 349.970 4.000 ;
    END
  END clk
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1049.350 0.000 1049.630 4.000 ;
    END
  END reset
  PIN rx
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 349.690 1396.000 349.970 1400.000 ;
    END
  END rx
  PIN tx
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1049.350 1396.000 1049.630 1400.000 ;
    END
  END tx
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 1387.440 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 1387.440 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 5.330 1383.065 1394.450 1385.895 ;
        RECT 5.330 1377.625 1394.450 1380.455 ;
        RECT 5.330 1372.185 1394.450 1375.015 ;
        RECT 5.330 1366.745 1394.450 1369.575 ;
        RECT 5.330 1361.305 1394.450 1364.135 ;
        RECT 5.330 1355.865 1394.450 1358.695 ;
        RECT 5.330 1350.425 1394.450 1353.255 ;
        RECT 5.330 1344.985 1394.450 1347.815 ;
        RECT 5.330 1339.545 1394.450 1342.375 ;
        RECT 5.330 1334.105 1394.450 1336.935 ;
        RECT 5.330 1328.665 1394.450 1331.495 ;
        RECT 5.330 1323.225 1394.450 1326.055 ;
        RECT 5.330 1317.785 1394.450 1320.615 ;
        RECT 5.330 1312.345 1394.450 1315.175 ;
        RECT 5.330 1306.905 1394.450 1309.735 ;
        RECT 5.330 1301.465 1394.450 1304.295 ;
        RECT 5.330 1296.025 1394.450 1298.855 ;
        RECT 5.330 1290.585 1394.450 1293.415 ;
        RECT 5.330 1285.145 1394.450 1287.975 ;
        RECT 5.330 1279.705 1394.450 1282.535 ;
        RECT 5.330 1274.265 1394.450 1277.095 ;
        RECT 5.330 1268.825 1394.450 1271.655 ;
        RECT 5.330 1263.385 1394.450 1266.215 ;
        RECT 5.330 1257.945 1394.450 1260.775 ;
        RECT 5.330 1252.505 1394.450 1255.335 ;
        RECT 5.330 1247.065 1394.450 1249.895 ;
        RECT 5.330 1241.625 1394.450 1244.455 ;
        RECT 5.330 1236.185 1394.450 1239.015 ;
        RECT 5.330 1230.745 1394.450 1233.575 ;
        RECT 5.330 1225.305 1394.450 1228.135 ;
        RECT 5.330 1219.865 1394.450 1222.695 ;
        RECT 5.330 1214.425 1394.450 1217.255 ;
        RECT 5.330 1208.985 1394.450 1211.815 ;
        RECT 5.330 1203.545 1394.450 1206.375 ;
        RECT 5.330 1198.105 1394.450 1200.935 ;
        RECT 5.330 1192.665 1394.450 1195.495 ;
        RECT 5.330 1187.225 1394.450 1190.055 ;
        RECT 5.330 1181.785 1394.450 1184.615 ;
        RECT 5.330 1176.345 1394.450 1179.175 ;
        RECT 5.330 1170.905 1394.450 1173.735 ;
        RECT 5.330 1165.465 1394.450 1168.295 ;
        RECT 5.330 1160.025 1394.450 1162.855 ;
        RECT 5.330 1154.585 1394.450 1157.415 ;
        RECT 5.330 1149.145 1394.450 1151.975 ;
        RECT 5.330 1143.705 1394.450 1146.535 ;
        RECT 5.330 1138.265 1394.450 1141.095 ;
        RECT 5.330 1132.825 1394.450 1135.655 ;
        RECT 5.330 1127.385 1394.450 1130.215 ;
        RECT 5.330 1121.945 1394.450 1124.775 ;
        RECT 5.330 1116.505 1394.450 1119.335 ;
        RECT 5.330 1111.065 1394.450 1113.895 ;
        RECT 5.330 1105.625 1394.450 1108.455 ;
        RECT 5.330 1100.185 1394.450 1103.015 ;
        RECT 5.330 1094.745 1394.450 1097.575 ;
        RECT 5.330 1089.305 1394.450 1092.135 ;
        RECT 5.330 1083.865 1394.450 1086.695 ;
        RECT 5.330 1078.425 1394.450 1081.255 ;
        RECT 5.330 1072.985 1394.450 1075.815 ;
        RECT 5.330 1067.545 1394.450 1070.375 ;
        RECT 5.330 1062.105 1394.450 1064.935 ;
        RECT 5.330 1056.665 1394.450 1059.495 ;
        RECT 5.330 1051.225 1394.450 1054.055 ;
        RECT 5.330 1045.785 1394.450 1048.615 ;
        RECT 5.330 1040.345 1394.450 1043.175 ;
        RECT 5.330 1034.905 1394.450 1037.735 ;
        RECT 5.330 1029.465 1394.450 1032.295 ;
        RECT 5.330 1024.025 1394.450 1026.855 ;
        RECT 5.330 1018.585 1394.450 1021.415 ;
        RECT 5.330 1013.145 1394.450 1015.975 ;
        RECT 5.330 1007.705 1394.450 1010.535 ;
        RECT 5.330 1002.265 1394.450 1005.095 ;
        RECT 5.330 996.825 1394.450 999.655 ;
        RECT 5.330 991.385 1394.450 994.215 ;
        RECT 5.330 985.945 1394.450 988.775 ;
        RECT 5.330 980.505 1394.450 983.335 ;
        RECT 5.330 975.065 1394.450 977.895 ;
        RECT 5.330 969.625 1394.450 972.455 ;
        RECT 5.330 964.185 1394.450 967.015 ;
        RECT 5.330 958.745 1394.450 961.575 ;
        RECT 5.330 953.305 1394.450 956.135 ;
        RECT 5.330 947.865 1394.450 950.695 ;
        RECT 5.330 942.425 1394.450 945.255 ;
        RECT 5.330 936.985 1394.450 939.815 ;
        RECT 5.330 931.545 1394.450 934.375 ;
        RECT 5.330 926.105 1394.450 928.935 ;
        RECT 5.330 920.665 1394.450 923.495 ;
        RECT 5.330 915.225 1394.450 918.055 ;
        RECT 5.330 909.785 1394.450 912.615 ;
        RECT 5.330 904.345 1394.450 907.175 ;
        RECT 5.330 898.905 1394.450 901.735 ;
        RECT 5.330 893.465 1394.450 896.295 ;
        RECT 5.330 888.025 1394.450 890.855 ;
        RECT 5.330 882.585 1394.450 885.415 ;
        RECT 5.330 877.145 1394.450 879.975 ;
        RECT 5.330 871.705 1394.450 874.535 ;
        RECT 5.330 866.265 1394.450 869.095 ;
        RECT 5.330 860.825 1394.450 863.655 ;
        RECT 5.330 855.385 1394.450 858.215 ;
        RECT 5.330 849.945 1394.450 852.775 ;
        RECT 5.330 844.505 1394.450 847.335 ;
        RECT 5.330 839.065 1394.450 841.895 ;
        RECT 5.330 833.625 1394.450 836.455 ;
        RECT 5.330 828.185 1394.450 831.015 ;
        RECT 5.330 822.745 1394.450 825.575 ;
        RECT 5.330 817.305 1394.450 820.135 ;
        RECT 5.330 811.865 1394.450 814.695 ;
        RECT 5.330 806.425 1394.450 809.255 ;
        RECT 5.330 800.985 1394.450 803.815 ;
        RECT 5.330 795.545 1394.450 798.375 ;
        RECT 5.330 790.105 1394.450 792.935 ;
        RECT 5.330 784.665 1394.450 787.495 ;
        RECT 5.330 779.225 1394.450 782.055 ;
        RECT 5.330 773.785 1394.450 776.615 ;
        RECT 5.330 768.345 1394.450 771.175 ;
        RECT 5.330 762.905 1394.450 765.735 ;
        RECT 5.330 757.465 1394.450 760.295 ;
        RECT 5.330 752.025 1394.450 754.855 ;
        RECT 5.330 746.585 1394.450 749.415 ;
        RECT 5.330 741.145 1394.450 743.975 ;
        RECT 5.330 735.705 1394.450 738.535 ;
        RECT 5.330 730.265 1394.450 733.095 ;
        RECT 5.330 724.825 1394.450 727.655 ;
        RECT 5.330 719.385 1394.450 722.215 ;
        RECT 5.330 713.945 1394.450 716.775 ;
        RECT 5.330 708.505 1394.450 711.335 ;
        RECT 5.330 703.065 1394.450 705.895 ;
        RECT 5.330 697.625 1394.450 700.455 ;
        RECT 5.330 692.185 1394.450 695.015 ;
        RECT 5.330 686.745 1394.450 689.575 ;
        RECT 5.330 681.305 1394.450 684.135 ;
        RECT 5.330 675.865 1394.450 678.695 ;
        RECT 5.330 670.425 1394.450 673.255 ;
        RECT 5.330 664.985 1394.450 667.815 ;
        RECT 5.330 659.545 1394.450 662.375 ;
        RECT 5.330 654.105 1394.450 656.935 ;
        RECT 5.330 648.665 1394.450 651.495 ;
        RECT 5.330 643.225 1394.450 646.055 ;
        RECT 5.330 637.785 1394.450 640.615 ;
        RECT 5.330 632.345 1394.450 635.175 ;
        RECT 5.330 626.905 1394.450 629.735 ;
        RECT 5.330 621.465 1394.450 624.295 ;
        RECT 5.330 616.025 1394.450 618.855 ;
        RECT 5.330 610.585 1394.450 613.415 ;
        RECT 5.330 605.145 1394.450 607.975 ;
        RECT 5.330 599.705 1394.450 602.535 ;
        RECT 5.330 594.265 1394.450 597.095 ;
        RECT 5.330 588.825 1394.450 591.655 ;
        RECT 5.330 583.385 1394.450 586.215 ;
        RECT 5.330 577.945 1394.450 580.775 ;
        RECT 5.330 572.505 1394.450 575.335 ;
        RECT 5.330 567.065 1394.450 569.895 ;
        RECT 5.330 561.625 1394.450 564.455 ;
        RECT 5.330 556.185 1394.450 559.015 ;
        RECT 5.330 550.745 1394.450 553.575 ;
        RECT 5.330 545.305 1394.450 548.135 ;
        RECT 5.330 539.865 1394.450 542.695 ;
        RECT 5.330 534.425 1394.450 537.255 ;
        RECT 5.330 528.985 1394.450 531.815 ;
        RECT 5.330 523.545 1394.450 526.375 ;
        RECT 5.330 518.105 1394.450 520.935 ;
        RECT 5.330 512.665 1394.450 515.495 ;
        RECT 5.330 507.225 1394.450 510.055 ;
        RECT 5.330 501.785 1394.450 504.615 ;
        RECT 5.330 496.345 1394.450 499.175 ;
        RECT 5.330 490.905 1394.450 493.735 ;
        RECT 5.330 485.465 1394.450 488.295 ;
        RECT 5.330 480.025 1394.450 482.855 ;
        RECT 5.330 474.585 1394.450 477.415 ;
        RECT 5.330 469.145 1394.450 471.975 ;
        RECT 5.330 463.705 1394.450 466.535 ;
        RECT 5.330 458.265 1394.450 461.095 ;
        RECT 5.330 452.825 1394.450 455.655 ;
        RECT 5.330 447.385 1394.450 450.215 ;
        RECT 5.330 441.945 1394.450 444.775 ;
        RECT 5.330 436.505 1394.450 439.335 ;
        RECT 5.330 431.065 1394.450 433.895 ;
        RECT 5.330 425.625 1394.450 428.455 ;
        RECT 5.330 420.185 1394.450 423.015 ;
        RECT 5.330 414.745 1394.450 417.575 ;
        RECT 5.330 409.305 1394.450 412.135 ;
        RECT 5.330 403.865 1394.450 406.695 ;
        RECT 5.330 398.425 1394.450 401.255 ;
        RECT 5.330 392.985 1394.450 395.815 ;
        RECT 5.330 387.545 1394.450 390.375 ;
        RECT 5.330 382.105 1394.450 384.935 ;
        RECT 5.330 376.665 1394.450 379.495 ;
        RECT 5.330 371.225 1394.450 374.055 ;
        RECT 5.330 365.785 1394.450 368.615 ;
        RECT 5.330 360.345 1394.450 363.175 ;
        RECT 5.330 354.905 1394.450 357.735 ;
        RECT 5.330 349.465 1394.450 352.295 ;
        RECT 5.330 344.025 1394.450 346.855 ;
        RECT 5.330 338.585 1394.450 341.415 ;
        RECT 5.330 333.145 1394.450 335.975 ;
        RECT 5.330 327.705 1394.450 330.535 ;
        RECT 5.330 322.265 1394.450 325.095 ;
        RECT 5.330 316.825 1394.450 319.655 ;
        RECT 5.330 311.385 1394.450 314.215 ;
        RECT 5.330 305.945 1394.450 308.775 ;
        RECT 5.330 300.505 1394.450 303.335 ;
        RECT 5.330 295.065 1394.450 297.895 ;
        RECT 5.330 289.625 1394.450 292.455 ;
        RECT 5.330 284.185 1394.450 287.015 ;
        RECT 5.330 278.745 1394.450 281.575 ;
        RECT 5.330 273.305 1394.450 276.135 ;
        RECT 5.330 267.865 1394.450 270.695 ;
        RECT 5.330 262.425 1394.450 265.255 ;
        RECT 5.330 256.985 1394.450 259.815 ;
        RECT 5.330 251.545 1394.450 254.375 ;
        RECT 5.330 246.105 1394.450 248.935 ;
        RECT 5.330 240.665 1394.450 243.495 ;
        RECT 5.330 235.225 1394.450 238.055 ;
        RECT 5.330 229.785 1394.450 232.615 ;
        RECT 5.330 224.345 1394.450 227.175 ;
        RECT 5.330 218.905 1394.450 221.735 ;
        RECT 5.330 213.465 1394.450 216.295 ;
        RECT 5.330 208.025 1394.450 210.855 ;
        RECT 5.330 202.585 1394.450 205.415 ;
        RECT 5.330 197.145 1394.450 199.975 ;
        RECT 5.330 191.705 1394.450 194.535 ;
        RECT 5.330 186.265 1394.450 189.095 ;
        RECT 5.330 180.825 1394.450 183.655 ;
        RECT 5.330 175.385 1394.450 178.215 ;
        RECT 5.330 169.945 1394.450 172.775 ;
        RECT 5.330 164.505 1394.450 167.335 ;
        RECT 5.330 159.065 1394.450 161.895 ;
        RECT 5.330 153.625 1394.450 156.455 ;
        RECT 5.330 148.185 1394.450 151.015 ;
        RECT 5.330 142.745 1394.450 145.575 ;
        RECT 5.330 137.305 1394.450 140.135 ;
        RECT 5.330 131.865 1394.450 134.695 ;
        RECT 5.330 126.425 1394.450 129.255 ;
        RECT 5.330 120.985 1394.450 123.815 ;
        RECT 5.330 115.545 1394.450 118.375 ;
        RECT 5.330 110.105 1394.450 112.935 ;
        RECT 5.330 104.665 1394.450 107.495 ;
        RECT 5.330 99.225 1394.450 102.055 ;
        RECT 5.330 93.785 1394.450 96.615 ;
        RECT 5.330 88.345 1394.450 91.175 ;
        RECT 5.330 82.905 1394.450 85.735 ;
        RECT 5.330 77.465 1394.450 80.295 ;
        RECT 5.330 72.025 1394.450 74.855 ;
        RECT 5.330 66.585 1394.450 69.415 ;
        RECT 5.330 61.145 1394.450 63.975 ;
        RECT 5.330 55.705 1394.450 58.535 ;
        RECT 5.330 50.265 1394.450 53.095 ;
        RECT 5.330 44.825 1394.450 47.655 ;
        RECT 5.330 39.385 1394.450 42.215 ;
        RECT 5.330 33.945 1394.450 36.775 ;
        RECT 5.330 28.505 1394.450 31.335 ;
        RECT 5.330 23.065 1394.450 25.895 ;
        RECT 5.330 17.625 1394.450 20.455 ;
        RECT 5.330 12.185 1394.450 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 1394.260 1387.285 ;
      LAYER met1 ;
        RECT 5.520 10.640 1394.260 1387.440 ;
      LAYER met2 ;
        RECT 9.300 1395.720 349.410 1396.000 ;
        RECT 350.250 1395.720 1049.070 1396.000 ;
        RECT 1049.910 1395.720 1390.020 1396.000 ;
        RECT 9.300 4.280 1390.020 1395.720 ;
        RECT 9.300 4.000 349.410 4.280 ;
        RECT 350.250 4.000 1049.070 4.280 ;
        RECT 1049.910 4.000 1390.020 4.280 ;
      LAYER met3 ;
        RECT 14.785 10.715 1384.995 1387.365 ;
      LAYER met4 ;
        RECT 94.135 11.735 97.440 1327.865 ;
        RECT 99.840 11.735 174.240 1327.865 ;
        RECT 176.640 11.735 251.040 1327.865 ;
        RECT 253.440 11.735 327.840 1327.865 ;
        RECT 330.240 11.735 404.640 1327.865 ;
        RECT 407.040 11.735 481.440 1327.865 ;
        RECT 483.840 11.735 558.240 1327.865 ;
        RECT 560.640 11.735 635.040 1327.865 ;
        RECT 637.440 11.735 711.840 1327.865 ;
        RECT 714.240 11.735 788.640 1327.865 ;
        RECT 791.040 11.735 865.440 1327.865 ;
        RECT 867.840 11.735 942.240 1327.865 ;
        RECT 944.640 11.735 1019.040 1327.865 ;
        RECT 1021.440 11.735 1095.840 1327.865 ;
        RECT 1098.240 11.735 1172.640 1327.865 ;
        RECT 1175.040 11.735 1249.440 1327.865 ;
        RECT 1251.840 11.735 1326.240 1327.865 ;
        RECT 1328.640 11.735 1378.785 1327.865 ;
  END
END leaf_chip
END LIBRARY

